module sobel3x3det(input [7:0] z1,
					input [7:0] z2,
					input [7:0] z3,
					input [7:0] z4,
					input [7:0] z5,
					input [7:0] z6,
					output [7:0] z_out
					);


	assign z_out = 8'b1;

endmodule